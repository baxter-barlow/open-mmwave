* PMIC behavioral model
VIN 1 0 DC 5
E3V3 2 0 1 0 0.66
E1V8 3 0 1 0 0.36
E1V2 4 0 1 0 0.24
E1V0 5 0 1 0 0.20
RLOAD3V3 2 0 33
RLOAD1V8 3 0 18
RLOAD1V2 4 0 12
RLOAD1V0 5 0 10
.op
.end
