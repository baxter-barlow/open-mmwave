* Power input ORing model
.include models/nsr20f30nxt5g.lib
VUSB 1 0 DC 5
VHD 2 0 DC 5
D1 1 3 NSR20F30NXT5G
D2 2 3 NSR20F30NXT5G
RLOAD 3 0 10
.op
.end
